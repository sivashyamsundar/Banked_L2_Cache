package L2manager;


